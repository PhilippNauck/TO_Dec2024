** sch_path: /ALL/Xschem/amps.xyce/hAMPsdiff_as1_3.5mA_15dB.sch
.subckt h_diff_15dB in VSS VDD sink ip op vGND
*.PININFO in:I VSS:B VDD:B sink:B ip:I op:O vGND:B
C1 net3 net2 10f
Q7 net2 in net7 net7 npn13G2 Nx=1
Q8 net3 ip net8 net8 npn13G2 Nx=1
R4 VDD net2 2e3
R5 VDD net3 2e3
R1 VDD net1 55e3
R2 vGND ip 10e3
R3 vGND in 10e3
R9 vGND VSS 20e3
R15 VDD vGND 20e3
Q9 net4 net1 VSS VSS npn13G2 Nx=1
Q5 net4 net1 VSS VSS npn13G2 Nx=1
Q3 VDD net2 net10 net10 npn13G2 Nx=1
Q4 VDD net3 net9 net9 npn13G2 Nx=1
Q10 net6 net5 VSS VSS npn13G2 Nx=1
Q11 op net6 VSS VSS npn13G2 Nx=6
Q12 net5 net5 VSS VSS npn13G2 Nx=1
R10 net7 net4 33
R12 net8 net4 33
R6 net10 net5 4e3
R8 net9 net6 4e3
Q1 net1 net1 VSS VSS npn13G2 Nx=1
R7 net10 net11 8e3
C2 net5 net11 .45e-15
**** begin user architecture code


**** end user architecture code
.ends
.end
